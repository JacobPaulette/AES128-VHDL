library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity mul9 is 
port(
	x: in std_logic_vector(7 downto 0);
	y: out std_logic_vector(7 downto 0)
); 
end mul9;

architecture mul9behavior of mul9 is
    subtype BYTE is std_logic_vector(7 downto 0);
    type LUT is array (0 to 255) of BYTE;
    constant mul9lut: LUT := (
"00000000","00001001","00010010","00011011","00100100","00101101","00110110","00111111",
"01001000","01000001","01011010","01010011","01101100","01100101","01111110","01110111",
"10010000","10011001","10000010","10001011","10110100","10111101","10100110","10101111",
"11011000","11010001","11001010","11000011","11111100","11110101","11101110","11100111",
"00111011","00110010","00101001","00100000","00011111","00010110","00001101","00000100",
"01110011","01111010","01100001","01101000","01010111","01011110","01000101","01001100",
"10101011","10100010","10111001","10110000","10001111","10000110","10011101","10010100",
"11100011","11101010","11110001","11111000","11000111","11001110","11010101","11011100",
"01110110","01111111","01100100","01101101","01010010","01011011","01000000","01001001",
"00111110","00110111","00101100","00100101","00011010","00010011","00001000","00000001",
"11100110","11101111","11110100","11111101","11000010","11001011","11010000","11011001",
"10101110","10100111","10111100","10110101","10001010","10000011","10011000","10010001",
"01001101","01000100","01011111","01010110","01101001","01100000","01111011","01110010",
"00000101","00001100","00010111","00011110","00100001","00101000","00110011","00111010",
"11011101","11010100","11001111","11000110","11111001","11110000","11101011","11100010",
"10010101","10011100","10000111","10001110","10110001","10111000","10100011","10101010",
"11101100","11100101","11111110","11110111","11001000","11000001","11011010","11010011",
"10100100","10101101","10110110","10111111","10000000","10001001","10010010","10011011",
"01111100","01110101","01101110","01100111","01011000","01010001","01001010","01000011",
"00110100","00111101","00100110","00101111","00010000","00011001","00000010","00001011",
"11010111","11011110","11000101","11001100","11110011","11111010","11100001","11101000",
"10011111","10010110","10001101","10000100","10111011","10110010","10101001","10100000",
"01000111","01001110","01010101","01011100","01100011","01101010","01110001","01111000",
"00001111","00000110","00011101","00010100","00101011","00100010","00111001","00110000",
"10011010","10010011","10001000","10000001","10111110","10110111","10101100","10100101",
"11010010","11011011","11000000","11001001","11110110","11111111","11100100","11101101",
"00001010","00000011","00011000","00010001","00101110","00100111","00111100","00110101",
"01000010","01001011","01010000","01011001","01100110","01101111","01110100","01111101",
"10100001","10101000","10110011","10111010","10000101","10001100","10010111","10011110",
"11101001","11100000","11111011","11110010","11001101","11000100","11011111","11010110",
"00110001","00111000","00100011","00101010","00010101","00011100","00000111","00001110",
"01111001","01110000","01101011","01100010","01011101","01010100","01001111","01000110"
);
begin
	y <= mul9lut(TO_INTEGER(unsigned(x)));
end;

