library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity mul13 is 
port(
	x: in std_logic_vector(7 downto 0);
	y: out std_logic_vector(7 downto 0)
); 
end mul13;

architecture mul13behavior of mul13 is
    subtype BYTE is std_logic_vector(7 downto 0);
    type LUT is array (0 to 255) of BYTE;
    constant mul13lut: LUT := (
"00000000","00001101","00011010","00010111","00110100","00111001","00101110","00100011",
"01101000","01100101","01110010","01111111","01011100","01010001","01000110","01001011",
"11010000","11011101","11001010","11000111","11100100","11101001","11111110","11110011",
"10111000","10110101","10100010","10101111","10001100","10000001","10010110","10011011",
"10111011","10110110","10100001","10101100","10001111","10000010","10010101","10011000",
"11010011","11011110","11001001","11000100","11100111","11101010","11111101","11110000",
"01101011","01100110","01110001","01111100","01011111","01010010","01000101","01001000",
"00000011","00001110","00011001","00010100","00110111","00111010","00101101","00100000",
"01101101","01100000","01110111","01111010","01011001","01010100","01000011","01001110",
"00000101","00001000","00011111","00010010","00110001","00111100","00101011","00100110",
"10111101","10110000","10100111","10101010","10001001","10000100","10010011","10011110",
"11010101","11011000","11001111","11000010","11100001","11101100","11111011","11110110",
"11010110","11011011","11001100","11000001","11100010","11101111","11111000","11110101",
"10111110","10110011","10100100","10101001","10001010","10000111","10010000","10011101",
"00000110","00001011","00011100","00010001","00110010","00111111","00101000","00100101",
"01101110","01100011","01110100","01111001","01011010","01010111","01000000","01001101",
"11011010","11010111","11000000","11001101","11101110","11100011","11110100","11111001",
"10110010","10111111","10101000","10100101","10000110","10001011","10011100","10010001",
"00001010","00000111","00010000","00011101","00111110","00110011","00100100","00101001",
"01100010","01101111","01111000","01110101","01010110","01011011","01001100","01000001",
"01100001","01101100","01111011","01110110","01010101","01011000","01001111","01000010",
"00001001","00000100","00010011","00011110","00111101","00110000","00100111","00101010",
"10110001","10111100","10101011","10100110","10000101","10001000","10011111","10010010",
"11011001","11010100","11000011","11001110","11101101","11100000","11110111","11111010",
"10110111","10111010","10101101","10100000","10000011","10001110","10011001","10010100",
"11011111","11010010","11000101","11001000","11101011","11100110","11110001","11111100",
"01100111","01101010","01111101","01110000","01010011","01011110","01001001","01000100",
"00001111","00000010","00010101","00011000","00111011","00110110","00100001","00101100",
"00001100","00000001","00010110","00011011","00111000","00110101","00100010","00101111",
"01100100","01101001","01111110","01110011","01010000","01011101","01001010","01000111",
"11011100","11010001","11000110","11001011","11101000","11100101","11110010","11111111",
"10110100","10111001","10101110","10100011","10000000","10001101","10011010","10010111"
);
begin
	y <= mul13lut(TO_INTEGER(unsigned(x)));
end;

