library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity mul11 is 
port(
	x: in std_logic_vector(7 downto 0);
	y: out std_logic_vector(7 downto 0)
); 
end mul11;

architecture mul11behavior of mul11 is
    subtype BYTE is std_logic_vector(7 downto 0);
    type LUT is array (0 to 255) of BYTE;
    constant mul11lut: LUT := (
"00000000","00001011","00010110","00011101","00101100","00100111","00111010","00110001",
"01011000","01010011","01001110","01000101","01110100","01111111","01100010","01101001",
"10110000","10111011","10100110","10101101","10011100","10010111","10001010","10000001",
"11101000","11100011","11111110","11110101","11000100","11001111","11010010","11011001",
"01111011","01110000","01101101","01100110","01010111","01011100","01000001","01001010",
"00100011","00101000","00110101","00111110","00001111","00000100","00011001","00010010",
"11001011","11000000","11011101","11010110","11100111","11101100","11110001","11111010",
"10010011","10011000","10000101","10001110","10111111","10110100","10101001","10100010",
"11110110","11111101","11100000","11101011","11011010","11010001","11001100","11000111",
"10101110","10100101","10111000","10110011","10000010","10001001","10010100","10011111",
"01000110","01001101","01010000","01011011","01101010","01100001","01111100","01110111",
"00011110","00010101","00001000","00000011","00110010","00111001","00100100","00101111",
"10001101","10000110","10011011","10010000","10100001","10101010","10110111","10111100",
"11010101","11011110","11000011","11001000","11111001","11110010","11101111","11100100",
"00111101","00110110","00101011","00100000","00010001","00011010","00000111","00001100",
"01100101","01101110","01110011","01111000","01001001","01000010","01011111","01010100",
"11110111","11111100","11100001","11101010","11011011","11010000","11001101","11000110",
"10101111","10100100","10111001","10110010","10000011","10001000","10010101","10011110",
"01000111","01001100","01010001","01011010","01101011","01100000","01111101","01110110",
"00011111","00010100","00001001","00000010","00110011","00111000","00100101","00101110",
"10001100","10000111","10011010","10010001","10100000","10101011","10110110","10111101",
"11010100","11011111","11000010","11001001","11111000","11110011","11101110","11100101",
"00111100","00110111","00101010","00100001","00010000","00011011","00000110","00001101",
"01100100","01101111","01110010","01111001","01001000","01000011","01011110","01010101",
"00000001","00001010","00010111","00011100","00101101","00100110","00111011","00110000",
"01011001","01010010","01001111","01000100","01110101","01111110","01100011","01101000",
"10110001","10111010","10100111","10101100","10011101","10010110","10001011","10000000",
"11101001","11100010","11111111","11110100","11000101","11001110","11010011","11011000",
"01111010","01110001","01101100","01100111","01010110","01011101","01000000","01001011",
"00100010","00101001","00110100","00111111","00001110","00000101","00011000","00010011",
"11001010","11000001","11011100","11010111","11100110","11101101","11110000","11111011",
"10010010","10011001","10000100","10001111","10111110","10110101","10101000","10100011",
);
begin
	y <= mul11lut(TO_INTEGER(unsigned(x)));
end;

