library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity mul14 is 
port(
	x: in std_logic_vector(7 downto 0);
	y: out std_logic_vector(7 downto 0)
); 
end mul14;

architecture mul14behavior of mul14 is
    subtype BYTE is std_logic_vector(7 downto 0);
    type LUT is array (0 to 255) of BYTE;
    constant mul14lut: LUT := (
"00000000","00001110","00011100","00010010","00111000","00110110","00100100","00101010",
"01110000","01111110","01101100","01100010","01001000","01000110","01010100","01011010",
"11100000","11101110","11111100","11110010","11011000","11010110","11000100","11001010",
"10010000","10011110","10001100","10000010","10101000","10100110","10110100","10111010",
"11011011","11010101","11000111","11001001","11100011","11101101","11111111","11110001",
"10101011","10100101","10110111","10111001","10010011","10011101","10001111","10000001",
"00111011","00110101","00100111","00101001","00000011","00001101","00011111","00010001",
"01001011","01000101","01010111","01011001","01110011","01111101","01101111","01100001",
"10101101","10100011","10110001","10111111","10010101","10011011","10001001","10000111",
"11011101","11010011","11000001","11001111","11100101","11101011","11111001","11110111",
"01001101","01000011","01010001","01011111","01110101","01111011","01101001","01100111",
"00111101","00110011","00100001","00101111","00000101","00001011","00011001","00010111",
"01110110","01111000","01101010","01100100","01001110","01000000","01010010","01011100",
"00000110","00001000","00011010","00010100","00111110","00110000","00100010","00101100",
"10010110","10011000","10001010","10000100","10101110","10100000","10110010","10111100",
"11100110","11101000","11111010","11110100","11011110","11010000","11000010","11001100",
"01000001","01001111","01011101","01010011","01111001","01110111","01100101","01101011",
"00110001","00111111","00101101","00100011","00001001","00000111","00010101","00011011",
"10100001","10101111","10111101","10110011","10011001","10010111","10000101","10001011",
"11010001","11011111","11001101","11000011","11101001","11100111","11110101","11111011",
"10011010","10010100","10000110","10001000","10100010","10101100","10111110","10110000",
"11101010","11100100","11110110","11111000","11010010","11011100","11001110","11000000",
"01111010","01110100","01100110","01101000","01000010","01001100","01011110","01010000",
"00001010","00000100","00010110","00011000","00110010","00111100","00101110","00100000",
"11101100","11100010","11110000","11111110","11010100","11011010","11001000","11000110",
"10011100","10010010","10000000","10001110","10100100","10101010","10111000","10110110",
"00001100","00000010","00010000","00011110","00110100","00111010","00101000","00100110",
"01111100","01110010","01100000","01101110","01000100","01001010","01011000","01010110",
"00110111","00111001","00101011","00100101","00001111","00000001","00010011","00011101",
"01000111","01001001","01011011","01010101","01111111","01110001","01100011","01101101",
"11010111","11011001","11001011","11000101","11101111","11100001","11110011","11111101",
"10100111","10101001","10111011","10110101","10011111","10010001","10000011","10001101"
);
begin
	y <= mul14lut(TO_INTEGER(unsigned(x)));
end;

