library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity mul2 is 
port(
	x: in std_logic_vector(7 downto 0);
	y: out std_logic_vector(7 downto 0)
); 
end mul2;

architecture mul2behavior of mul2 is
    subtype BYTE is std_logic_vector(7 downto 0);
    type LUT is array (0 to 255) of BYTE;
    constant mul2lut: LUT := (
"00000000","00000010","00000100","00000110","00001000","00001010","00001100","00001110",
"00010000","00010010","00010100","00010110","00011000","00011010","00011100","00011110",
"00100000","00100010","00100100","00100110","00101000","00101010","00101100","00101110",
"00110000","00110010","00110100","00110110","00111000","00111010","00111100","00111110",
"01000000","01000010","01000100","01000110","01001000","01001010","01001100","01001110",
"01010000","01010010","01010100","01010110","01011000","01011010","01011100","01011110",
"01100000","01100010","01100100","01100110","01101000","01101010","01101100","01101110",
"01110000","01110010","01110100","01110110","01111000","01111010","01111100","01111110",
"10000000","10000010","10000100","10000110","10001000","10001010","10001100","10001110",
"10010000","10010010","10010100","10010110","10011000","10011010","10011100","10011110",
"10100000","10100010","10100100","10100110","10101000","10101010","10101100","10101110",
"10110000","10110010","10110100","10110110","10111000","10111010","10111100","10111110",
"11000000","11000010","11000100","11000110","11001000","11001010","11001100","11001110",
"11010000","11010010","11010100","11010110","11011000","11011010","11011100","11011110",
"11100000","11100010","11100100","11100110","11101000","11101010","11101100","11101110",
"11110000","11110010","11110100","11110110","11111000","11111010","11111100","11111110",
"00011011","00011001","00011111","00011101","00010011","00010001","00010111","00010101",
"00001011","00001001","00001111","00001101","00000011","00000001","00000111","00000101",
"00111011","00111001","00111111","00111101","00110011","00110001","00110111","00110101",
"00101011","00101001","00101111","00101101","00100011","00100001","00100111","00100101",
"01011011","01011001","01011111","01011101","01010011","01010001","01010111","01010101",
"01001011","01001001","01001111","01001101","01000011","01000001","01000111","01000101",
"01111011","01111001","01111111","01111101","01110011","01110001","01110111","01110101",
"01101011","01101001","01101111","01101101","01100011","01100001","01100111","01100101",
"10011011","10011001","10011111","10011101","10010011","10010001","10010111","10010101",
"10001011","10001001","10001111","10001101","10000011","10000001","10000111","10000101",
"10111011","10111001","10111111","10111101","10110011","10110001","10110111","10110101",
"10101011","10101001","10101111","10101101","10100011","10100001","10100111","10100101",
"11011011","11011001","11011111","11011101","11010011","11010001","11010111","11010101",
"11001011","11001001","11001111","11001101","11000011","11000001","11000111","11000101",
"11111011","11111001","11111111","11111101","11110011","11110001","11110111","11110101",
"11101011","11101001","11101111","11101101","11100011","11100001","11100111","11100101"
);

begin
	y <= mul2lut(TO_INTEGER(unsigned(x)));
end;

