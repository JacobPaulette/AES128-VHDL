library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity mul2 is 
port(
	x: in std_logic_vector(7 downto 0);
	y: out std_logic_vector(7 downto 0)
); 
end mul2;

architecture mul2behavior of mul2 is
    subtype BYTE is std_logic_vector(7 downto 0);
    type LUT is array (0 to 255) of BYTE;
    constant mul2lut: LUT := (
"00000000","00000011","00000110","00000101","00001100","00001111","00001010","00001001",
"00011000","00011011","00011110","00011101","00010100","00010111","00010010","00010001",
"00110000","00110011","00110110","00110101","00111100","00111111","00111010","00111001",
"00101000","00101011","00101110","00101101","00100100","00100111","00100010","00100001",
"01100000","01100011","01100110","01100101","01101100","01101111","01101010","01101001",
"01111000","01111011","01111110","01111101","01110100","01110111","01110010","01110001",
"01010000","01010011","01010110","01010101","01011100","01011111","01011010","01011001",
"01001000","01001011","01001110","01001101","01000100","01000111","01000010","01000001",
"11000000","11000011","11000110","11000101","11001100","11001111","11001010","11001001",
"11011000","11011011","11011110","11011101","11010100","11010111","11010010","11010001",
"11110000","11110011","11110110","11110101","11111100","11111111","11111010","11111001",
"11101000","11101011","11101110","11101101","11100100","11100111","11100010","11100001",
"10100000","10100011","10100110","10100101","10101100","10101111","10101010","10101001",
"10111000","10111011","10111110","10111101","10110100","10110111","10110010","10110001",
"10010000","10010011","10010110","10010101","10011100","10011111","10011010","10011001",
"10001000","10001011","10001110","10001101","10000100","10000111","10000010","10000001",
"10011011","10011000","10011101","10011110","10010111","10010100","10010001","10010010",
"10000011","10000000","10000101","10000110","10001111","10001100","10001001","10001010",
"10101011","10101000","10101101","10101110","10100111","10100100","10100001","10100010",
"10110011","10110000","10110101","10110110","10111111","10111100","10111001","10111010",
"11111011","11111000","11111101","11111110","11110111","11110100","11110001","11110010",
"11100011","11100000","11100101","11100110","11101111","11101100","11101001","11101010",
"11001011","11001000","11001101","11001110","11000111","11000100","11000001","11000010",
"11010011","11010000","11010101","11010110","11011111","11011100","11011001","11011010",
"01011011","01011000","01011101","01011110","01010111","01010100","01010001","01010010",
"01000011","01000000","01000101","01000110","01001111","01001100","01001001","01001010",
"01101011","01101000","01101101","01101110","01100111","01100100","01100001","01100010",
"01110011","01110000","01110101","01110110","01111111","01111100","01111001","01111010",
"00111011","00111000","00111101","00111110","00110111","00110100","00110001","00110010",
"00100011","00100000","00100101","00100110","00101111","00101100","00101001","00101010",
"00001011","00001000","00001101","00001110","00000111","00000100","00000001","00000010",
"00010011","00010000","00010101","00010110","00011111","00011100","00011001","00011010"
);
begin
	y <= mul2lut(TO_INTEGER(unsigned(x)));
end;

